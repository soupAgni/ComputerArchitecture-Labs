library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mux_4to1 is
    generic(N : integer := 32);
    Port ( SEL : in  STD_LOGIC_VECTOR (1 downto 0);
           A   : in  STD_LOGIC;
           B   : in  STD_LOGIC;
           C   : in  STD_LOGIC;
           D   : in  STD_LOGIC;
           X   : out STD_LOGIC);
end mux_4to1;

architecture Behavioral of mux_4to1 is
begin
   
   x <= A when SEL = "00" else
        B when SEL = "01" else
        C when SEL = "10" else
        D when SEL = "11" else
        '0';
   
end Behavioral;