use work.all;
library IEEE;
use IEEE.std_logic_1164.all;


entity multiplexer_c is
  
  generic(N : integer := 32);
  port(x         : in std_logic_vector(N-1 downto 0);
       A         : in std_logic_vector(N-1 downto 0);
       B         : in std_logic_vector(N-1 downto 0);
       Y         : out std_logic_vector(N-1 downto 0));

end multiplexer_c;

architecture dataflow of multiplexer_c is
  component multiplexer is
  
  port(x         : in std_logic;
       A         : in std_logic;
       B         : in std_logic;
       Y         : out std_logic);

end component;


  
begin

G1: for i in 0 to N-1 generate
  
  multiplexer_1 : multiplexer
  
  port map(
  
  x  => x(i),
  A  => A(i),
  B  => B(i),
  Y  => Y(i));
 
end generate;
  
end dataflow;
