use work.all;
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ALU_1bit_P2 is
    generic(N : integer := 1);
    Port ( A        : in  STD_LOGIC;
           B        : in  STD_LOGIC;
           Less     : in  STD_LOGIC;
           Cin      : in  STD_LOGIC;
           Op       : in  STD_LOGIC_VECTOR (2 downto 0);
           Ainvert  : in  STD_LOGIC;
           Binvert  : in  STD_LOGIC;
           Overflow : out STD_LOGIC;
           Set      : out STD_LOGIC;
           Result   : out STD_LOGIC;
           Carry_out:  out STD_LOGIC);
end ALU_1bit_P2;
---------------------------
architecture dataflow of ALU_1bit_P2 is
----------------------------  
  component multiplexer 
     port(x         : in std_logic;
       A         : in std_logic;
       B         : in std_logic;
       Y         : out std_logic);

  end component;
---------------------------  
  component or2 
  port(i_A          : in std_logic;
       i_B          : in std_logic;
       o_F          : out std_logic);

  end component;
----------------------------  
  component inv 
  port(i_A          : in std_logic;
       o_F          : out std_logic);
  end component;
----------------------------
  component and2
  port(i_A          : in std_logic;
       i_B          : in std_logic;
       o_F          : out std_logic);
  end component;
---------------------------
  component xor2 is

  port(i_A          : in std_logic;
       i_B          : in std_logic;
       o_F          : out std_logic);

  end component;
----------------------------
  COMPONENT mux_5to1_top 
    generic(N : integer := 1);
    Port ( SEL : in  STD_LOGIC_VECTOR (2 downto 0);
           A   : in  STD_LOGIC;
           B   : in  STD_LOGIC;
           C   : in  STD_LOGIC;
           D   : in  STD_LOGIC;
           E   : in  STD_LOGIC;
           X   : out STD_LOGIC);
end component;
 --------------------------- 
  component fullAdder_b 
  port(C_in      : in std_logic;
       A         : in std_logic;
       B         : in std_logic;
       C_out     : out std_logic;
       S_out     : out std_logic);
  end component;
 ----------------------------- 
  signal s_inv1, s_inv2, s_Ainv,s_Binv, s_And1, s_Or1, s_Adder, s_XOR, s_5to1mux: STD_LOGIC;
  signal temp : STD_LOGIC:= '0';
 ----------------------------- 
  begin 
    
    xor1 : xor2 
    port map(i_A   => A,
             i_B   => B,
             o_F   => s_XOR);
    
    inv1 : inv
    port map(i_A   => A,
             o_F   => s_inv1);
            
            
    inv2 : inv
    port map(i_A   => B,
             o_F   => s_inv2);
    
    mux1 :    multiplexer      
    port map( X => Ainvert,
              A   => A,
              B   => s_inv1,
              Y   => s_Ainv);   
              
    mux2 :   multiplexer       
    port map( X => Binvert,
              A   => B,
              B   => s_inv2,
              Y   => s_Binv);     
    
    and1 :   and2      
    port map(i_A  => s_Ainv,
             i_B  => s_Binv,
             o_F  => s_And1);
    or1 : or2        
    port map(i_A  => s_Ainv,
             i_B  => s_Binv,
             o_F  => s_Or1);
     
    fullAdder :   fullAdder_b
    port map(C_in  => Cin,
             A     => s_Ainv,
             B     => s_Binv,
             C_out => temp, 
             S_out => s_Adder);
             
    mux5to1 :  mux_5to1_top   
    port map( SEL => Op,
              A   => s_And1,
              B   => s_Or1,
              C   => s_Adder,
              D  =>  Less,
              E  =>  s_XOR,
              X   => s_5to1mux);
              
    Result <= s_5to1mux;          
    Set <= s_Adder;
    Overflow <= (s_Ainv and s_Binv and (not s_Adder)) or ((not s_Ainv) and (not s_Binv) and s_Adder);
    Carry_out <= temp;
      
end dataflow;